----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 2018/11/24 10:55:57
-- Design Name: 
-- Module Name: solve - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.std_logic_signed.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity display_test is port(
    ans : in std_logic_vector(8 downto 0);
    clk, flag, do : in std_logic;
    en: out std_logic_vector(5 downto 0);
    seg : out std_logic_vector(7 downto 0));
end display_test;

architecture behavioral of display_test is
    signal div_cnt: integer range 0 to 150 := 0;
    signal div_clk: std_logic := '0';
    signal seg1, seg2, seg3, seg4, seg5, seg6: std_logic_vector(7 downto 0);
    signal disp_bit : std_logic_vector(3 downto 0) := "0000";
    signal new_bit : std_logic_vector(3 downto 0);
begin
    process (clk)
    begin
        if clk'event and clk = '1' then
           if div_cnt = 100 then
                    div_clk <= not div_clk;
                    div_cnt <= 0;
           else 
                    div_cnt <= div_cnt + 1;
           end if;
       end if;
    end process;
    
    seg1 <= "01000000" when flag = '1' else "00000000";
    seg2 <= "10000110" when ans(6) = '1' else "10111111";
    
    process(ans)
    begin
        case ans(5 downto 0) is
            when "000000" =>
                seg3 <= "00111111";
                seg4 <= "00111111";
                seg5 <= "00111111";
                seg6 <= "00111111"; --0.0000
            when "000001" =>
                seg3 <= "00111111";
                seg4 <= "00000110";
                seg5 <= "01101101";
                seg6 <= "01111101"; --0.0156 
            when "000010" =>
                seg3 <= "00111111";
                seg4 <= "01001111";
                seg5 <= "00000110";
                seg6 <= "01011011"; --0.0312
            when "000011" =>
                seg3 <= "00111111";
                seg4 <= "01100110";
                seg5 <= "01111101";
                seg6 <= "01111111"; --0.0468    
            when "000100" =>
                seg3 <= "00111111";
                seg4 <= "01111101";
                seg5 <= "01011011";
                seg6 <= "01101101"; --0.0625
            when "000101" =>
                seg3 <= "00111111";
                seg4 <= "00000111";
                seg5 <= "01111111";
                seg6 <= "00000110"; --0.0781
            when "000110" =>
                seg3 <= "00111111";
                seg4 <= "01101111";
                seg5 <= "01001111";
                seg6 <= "00000111"; --0.0937
            when "000111" =>
                seg3 <= "00000110";
                seg4 <= "00111111";
                seg5 <= "01101111";
                seg6 <= "01001111"; --0.1093
           when "001000" =>
                seg3 <= "00000110";
                seg4 <= "01011011";
                seg5 <= "01101101";
                seg6 <= "00111111"; --0.1250
           when "001001" =>
                seg3 <= "00000110";
                seg4 <= "01100110";
                seg5 <= "00111111";
                seg6 <= "01111101"; --0.1406
           when "001010" =>
                seg3 <= "00000110";
                seg4 <= "01101101";
                seg5 <= "01111101";
                seg6 <= "01011011"; --0.1562
           when "001011" =>
                seg3 <= "00000110";
                seg4 <= "00000111";
                seg5 <= "00000110";
                seg6 <= "01111111"; --0.1718
           when "001100" =>
                seg3 <= "00000110";
                seg4 <= "01111111";
                seg5 <= "00000111";
                seg6 <= "01101101"; --0.1875
           when "001101" =>
                seg3 <= "01011011";
                seg4 <= "00111111";
                seg5 <= "01001111";
                seg6 <= "00000110"; --0.2031
           when "001110" =>
                seg3 <= "01011011";
                seg4 <= "00000110";
                seg5 <= "01111111";
                seg6 <= "00000111"; --0.2187
          when "001111" =>
                seg3 <= "01011011";
                seg4 <= "01001111";
                seg5 <= "01100110";
                seg6 <= "01001111"; --0.2343
          when "010000" =>
                seg3 <= "01011011";
                seg4 <= "01101101";
                seg5 <= "00111111";
                seg6 <= "00111111"; --0.2500
          when "010001" =>
                seg3 <= "01011011";
                seg4 <= "01111101";
                seg5 <= "01101101";
                seg6 <= "01111101"; --0.2656
          when "010010" =>
                seg3 <= "01011011";
                seg4 <= "01111111";
                seg5 <= "00000110";
                seg6 <= "01011011"; --0.2812
          when "010011" =>
                seg3 <= "01011011";
                seg4 <= "01101111";
                seg5 <= "01111101";
                seg6 <= "01111111"; --0.2968
          when "010100" =>
                seg3 <= "01001111";
                seg4 <= "00000110";
                seg5 <= "01011011";
                seg6 <= "01101101"; --0.3125
          when "010101" =>
                seg3 <= "01001111";
                seg4 <= "01011011";
                seg5 <= "01111111";
                seg6 <= "00000110"; --0.3281
         when "010110" =>
                seg3 <= "01001111";
                seg4 <= "01100110";
                seg5 <= "01001111";
                seg6 <= "00000111"; --0.3437
         when "010111" =>
                seg3 <= "01001111";
                seg4 <= "01101101";
                seg5 <= "01101111";
                seg6 <= "01001111"; --0.3593
         when "011000" =>
                seg3 <= "01001111";
                seg4 <= "00000111";
                seg5 <= "01101101";
                seg6 <= "00111111"; --0.3750
         when "011001" =>
                seg3 <= "01001111";
                seg4 <= "01101111";
                seg5 <= "00111111";
                seg6 <= "01111101"; --0.3906
         when "011010" =>
                seg3 <= "01100110";
                seg4 <= "00111111";
                seg5 <= "01111101";
                seg6 <= "01011011"; --0.4062
         when "011011" =>
                seg3 <= "01100110";
                seg4 <= "01011011";
                seg5 <= "00000110";
                seg6 <= "01111111"; --0.4218
         when "011100" =>
                seg3 <= "01100110";
                seg4 <= "01001111";
                seg5 <= "00000111";
                seg6 <= "01101101"; --0.4375
         when "011101" =>
                seg3 <= "01100110";
                seg4 <= "01101101";
                seg5 <= "01001111";
                seg6 <= "00000110"; --0.4531
         when "011110" =>
                seg3 <= "01100110";
                seg4 <= "01111101";
                seg5 <= "01111111";
                seg6 <= "00000111"; --0.4687
         when "011111" =>
                seg3 <= "01100110";
                seg4 <= "01111111";
                seg5 <= "01100110";
                seg6 <= "01001111"; --0.4843
         when "100000" =>
                seg3 <= "01101101";
                seg4 <= "00111111";
                seg5 <= "00111111";
                seg6 <= "00111111"; --0.5000
            when "100001" =>
                seg3 <= "01101101";
                seg4 <= "00000110";
                seg5 <= "01101101";
                seg6 <= "01111101"; --0.5156 
            when "100010" =>
                seg3 <= "01101101";
                seg4 <= "01001111";
                seg5 <= "00000110";
                seg6 <= "01011011"; --0.5312
            when "100011" =>
                seg3 <= "01101101";
                seg4 <= "01100110";
                seg5 <= "01111101";
                seg6 <= "01111111"; --0.5468    
            when "100100" =>
                seg3 <= "01101101";
                seg4 <= "01111101";
                seg5 <= "01011011";
                seg6 <= "01101101"; --0.5625
            when "100101" =>
                seg3 <= "01101101";
                seg4 <= "00000111";
                seg5 <= "01111111";
                seg6 <= "00000110"; --0.5781
            when "100110" =>
                seg3 <= "01101101";
                seg4 <= "01101111";
                seg5 <= "01001111";
                seg6 <= "00000111"; --0.5937
            when "100111" =>
                seg3 <= "01111101";
                seg4 <= "00111111";
                seg5 <= "01101111";
                seg6 <= "01001111"; --0.6093
           when "101000" =>
                seg3 <= "01111101";
                seg4 <= "01011011";
                seg5 <= "01101101";
                seg6 <= "00111111"; --0.6250
           when "101001" =>
                seg3 <= "01111101";
                seg4 <= "01100110";
                seg5 <= "00111111";
                seg6 <= "01111101"; --0.6406
           when "101010" =>
                seg3 <= "01111101";
                seg4 <= "01101101";
                seg5 <= "01111101";
                seg6 <= "01011011"; --0.6562
           when "101011" =>
                seg3 <= "01111101";
                seg4 <= "00000111";
                seg5 <= "00000110";
                seg6 <= "01111111"; --0.6718
           when "101100" =>
                seg3 <= "01111101";
                seg4 <= "01111111";
                seg5 <= "00000111";
                seg6 <= "01101101"; --0.6875
           when "101101" =>
                seg3 <= "00000111";
                seg4 <= "00111111";
                seg5 <= "01001111";
                seg6 <= "00000110"; --0.7031
           when "101110" =>
                seg3 <= "00000111";
                seg4 <= "00000110";
                seg5 <= "01111111";
                seg6 <= "00000111"; --0.7187
          when "101111" =>
                seg3 <= "00000111";
                seg4 <= "01001111";
                seg5 <= "01100110";
                seg6 <= "01001111"; --0.7343
          when "110000" =>
                seg3 <= "00000111";
                seg4 <= "01101101";
                seg5 <= "00111111";
                seg6 <= "00111111"; --0.7500
          when "110001" =>
                seg3 <= "00000111";
                seg4 <= "01111101";
                seg5 <= "01101101";
                seg6 <= "01111101"; --0.7656
          when "110010" =>
                seg3 <= "00000111";
                seg4 <= "01111111";
                seg5 <= "00000110";
                seg6 <= "01011011"; --0.7812
          when "110011" =>
                seg3 <= "00000111";
                seg4 <= "01101111";
                seg5 <= "01111101";
                seg6 <= "01111111"; --0.7968
          when "110100" =>
                seg3 <= "01111111";
                seg4 <= "00000110";
                seg5 <= "01011011";
                seg6 <= "01101101"; --0.8125
          when "110101" =>
                seg3 <= "01111111";
                seg4 <= "01011011";
                seg5 <= "01111111";
                seg6 <= "00000110"; --0.8281
         when "110110" =>
                seg3 <= "01111111";
                seg4 <= "01100110";
                seg5 <= "01001111";
                seg6 <= "00000111"; --0.8437
         when "110111" =>
                seg3 <= "01111111";
                seg4 <= "01101101";
                seg5 <= "01101111";
                seg6 <= "01001111"; --0.8593
         when "111000" =>
                seg3 <= "01111111";
                seg4 <= "00000111";
                seg5 <= "01101101";
                seg6 <= "00111111"; --0.8750
         when "111001" =>
                seg3 <= "01111111";
                seg4 <= "01101111";
                seg5 <= "00111111";
                seg6 <= "01111101"; --0.8906
         when "111010" =>
                seg3 <= "01101111";
                seg4 <= "00111111";
                seg5 <= "01111101";
                seg6 <= "01011011"; --0.9062
         when "111011" =>
                seg3 <= "01101111";
                seg4 <= "01011011";
                seg5 <= "00000110";
                seg6 <= "01111111"; --0.9218
         when "111100" =>
                seg3 <= "01101111";
                seg4 <= "01001111";
                seg5 <= "00000111";
                seg6 <= "01101101"; --0.9375
         when "111101" =>
                seg3 <= "01101111";
                seg4 <= "01101101";
                seg5 <= "01001111";
                seg6 <= "00000110"; --0.9531
         when "111110" =>
                seg3 <= "01101111";
                seg4 <= "01111101";
                seg5 <= "01111111";
                seg6 <= "00000111"; --0.9687
         when "111111" =>
                seg3 <= "01101111";
                seg4 <= "01111111";
                seg5 <= "01100110";
                seg6 <= "01001111"; --0.9843
         when others =>
                seg3 <= "00111111";
                seg4 <= "00111111";
                seg5 <= "00111111";
                seg6 <= "00111111";
        end case;
    end process;
    
    process(div_clk)
    begin
        if div_clk'event and div_clk = '1' then
            if do = '0' then
                disp_bit <= "0000";
            else
                case disp_bit is
                    when "0000" =>
                        en <= "111111";
                        seg <= "00000000";
                        new_bit <= disp_bit + '1';
                    when "0001" =>
                        en <= "111110";
                        new_bit <= disp_bit + '1';
                        seg <= seg6;
                    when "0010" =>
                        en <= "111101";
                        seg <= seg5;
                        new_bit <= disp_bit + '1';
                    when "0011" =>
                        en <= "111011";
                        seg <= seg4;
                        new_bit <= disp_bit + '1';
                    when "0100" =>
                        en <= "110111";
                        seg <= seg3;
                        new_bit <= disp_bit + '1';
                    when "0101" =>
                        en <= "101111";
                        seg <= seg2;
                        new_bit <= disp_bit + '1';
                    when "0110" =>
                        en <= "011111";
                        seg <= seg1;
                        new_bit <= "0001";
                    when others =>
                        en <= "111111"; 
                        seg <= "00000000";
                end case;  
                disp_bit <= new_bit;
            end if; 
        end if;
    end process;

end behavioral;